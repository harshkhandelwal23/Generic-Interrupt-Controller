package pkg;
  `include "uvm_macros.svh"
  import uvm_pkg::*;
  `include "../SEQ_LIB/interrupt_seq_item.sv"
  `include "../SEQ_LIB/interrupt_seq.sv"
  `include "reg_block.sv"
  `include "../SEQ_LIB/reg_seq_item.sv"
  `include "reg_adapter.sv"
  `include "../SEQ_LIB/reg_seq.sv"
  `include "reg_seqr.sv"
  `include "reg_driver.sv"
  `include "reg_monitor.sv"
  `include "reg_agent.sv"
  `include "interrupt_seqr.sv"
  `include "interrupt_driver.sv"
  `include "interrupt_monitor.sv"
  `include "int_out_monitor.sv"
  `include "interrupt_agent.sv"
  `include "int_out_agent.sv"
  `include "intc_scoreboard.sv"
  `include "interrupt_env.sv"
  `include "../SEQ_LIB/sanity_seq.sv"
  `include "../TEST/sanity_test.sv"
  `include "../TEST/reg_test.sv"
endpackage
