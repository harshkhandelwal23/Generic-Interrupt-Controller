`define no_of_sources 10
