`define no_of_sources 11
